../functional/vhdl.vhd